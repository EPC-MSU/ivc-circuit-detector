* Qucs 2.1.0 C:/dev/ivc-circuit-detector/circuit_classes/CR/CR.sch
.INCLUDE "C:/Program Files (x86)/Qucs-S/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
* Qucs 2.1.0  C:/dev/ivc-circuit-detector/circuit_classes/CR/CR.sch
C1 input 0  1N 
R1 input 0  1K
.control
set filetype=ascii
op
print all > spice4qucs.cir.dc_op
destroy all
quit
.endc
.end
