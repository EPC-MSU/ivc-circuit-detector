* Qucs 2.1.0 C:/dev/ivc-circuit-detector/circuit_classes/R_C/R_C.sch
.INCLUDE "C:/Program Files (x86)/Qucs-S/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
* Qucs 2.1.0  C:/dev/ivc-circuit-detector/circuit_classes/R_C/R_C.sch
R1 input _net0  1K
C1 0 _net0  1N 
.control
set filetype=ascii
op
print all > spice4qucs.cir.dc_op
destroy all
quit
.endc
.end
