* Qucs 25.2.0  C:/Users/volkov_pa/Desktop/workdir/ivc-circuit-detector/circuit_classes/D_C/D_C.sch
.INCLUDE "C:/Program Files/Qucs-S/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
C1 0 _net0  1N 
D1 input _net0 DMOD_D1 AREA=1.0
.MODEL DMOD_D1 D (Is=222P N=1.65 Cj0=0P M=0.0 Vj=0.7 Fc=0.5 Rs=68.6M Tt=5.76N Kf=0 Af=1 Bv=75 Ibv=1U Xti=3.0 Eg=1.11 Tcv=0.0 Trs=0.0 Ttt1=0.0 Ttt2=0.0 Tm1=0.0 Tm2=0.0 Tnom=26.85 )

.control

op
print v(input)   > spice4qucs.dc1.ngspice.dc.print
destroy all
reset

exit
.endc
.END
