* Qucs 2.1.0 C:/dev/ivc-circuit-detector/circuit_classes/DD_R_1N4148/DD_R_1N4148.sch
.INCLUDE "C:/Program Files (x86)/Qucs-S/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
* Qucs 2.1.0  C:/dev/ivc-circuit-detector/circuit_classes/DD_R_1N4148/DD_R_1N4148.sch
D_1N4148_1 _net0 input DMOD_D_1N4148_1 AREA=1.0 Temp=26.85
.MODEL DMOD_D_1N4148_1 D (Is=2.22e-10 N=1.65 Cj0=4e-12 M=0.333 Vj=0.7 Fc=0.5 Rs=0.0686 Tt=5.76e-09 Kf=0 Af=1 Bv=75 Ibv=1e-06 Xti=3 Eg=1.11 Tcv=0 Trs=0 Ttt1=0 Ttt2=0 Tm1=0 Tm2=0 Tnom=26.85 )
R1 0 _net0  1K
D_1N4148_2 input _net0 DMOD_D_1N4148_2 AREA=1.0 Temp=26.85
.MODEL DMOD_D_1N4148_2 D (Is=2.22e-10 N=1.65 Cj0=4e-12 M=0.333 Vj=0.7 Fc=0.5 Rs=0.0686 Tt=5.76e-09 Kf=0 Af=1 Bv=75 Ibv=1e-06 Xti=3 Eg=1.11 Tcv=0 Trs=0 Ttt1=0 Ttt2=0 Tm1=0 Tm2=0 Tnom=26.85 )
.control
set filetype=ascii
op
print all > spice4qucs.cir.dc_op
destroy all
quit
.endc
.end
